library verilog;
use verilog.vl_types.all;
entity half_adder_testbench is
end half_adder_testbench;
